*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'mhao' on Mon Oct 24 2016 at 18:47:37

*
* Globals.
*
.global VDD GROUND

*
* Component pathname : $UpdatedFiles/default.group/logic.views/AND
*
.subckt AND  OUT A B

        M1 OUT N$4 GROUND GROUND N L=.4u W=1.2u M=1
        M3 N$6 A GROUND GROUND N L=.4u W=2.4u M=1
        M5 N$4 B N$6 GROUND N L=.4u W=2.4u M=1
        M4 N$4 B VDD VDD P L=.4u W=2.4u M=1
        M6 N$4 A VDD VDD P L=.4u W=2.4u M=1
        M2 OUT N$4 VDD VDD P L=.4u W=2.4u M=1
.ends AND

*
* Component pathname : $UpdatedFiles/default.group/logic.views/inverter
*
.subckt INVERTER  OUT IN

        M2 OUT IN VDD VDD P L=0.4u W=3.6u M=1
        M1 OUT IN GROUND GROUND N L=0.4u W=1.2u M=1
.ends INVERTER

*
* Component pathname : $UpdatedFiles/default.group/logic.views/153_XOR
*
.subckt 153_XOR  XOR A B

        X_INVERTER1 XOR N$3 INVERTER
        M2 B A N$3 GROUND N L=0.4u W=1.2u M=2
        M4 A B N$3 GROUND N L=0.4u W=1.2u M=2
        M3 N$3 B N$2 VDD P L=0.4u W=2.4u M=2
        M1 N$2 A VDD VDD P L=0.4u W=2.4u M=2
.ends 153_XOR

*
* Component pathname : $UpdatedFiles/default.group/logic.views/Half-Adder
*
.subckt HALF-ADDER  C S X Y

        X_AND1 C Y X AND
        X_153_XOR1 S Y X 153_XOR
.ends HALF-ADDER

*
* Component pathname : $UpdatedFiles/default.group/logic.views/OR
*
.subckt OR  OUT A B

        M3 N$12 A GROUND GROUND N L=.4u W=1.2u M=1
        M1 N$12 B GROUND GROUND N L=.4u W=1.2u M=1
        M6 OUT N$12 VDD VDD P L=.4u W=2.4u M=1
        M5 OUT N$12 GROUND GROUND N L=.4u W=1.2u M=1
        M4 N$12 B N$8 VDD P L=.4u W=4.8u M=1
        M2 N$8 A VDD VDD P L=.4u W=4.8u M=1
.ends OR

*
* Component pathname : $UpdatedFiles/default.group/logic.views/Full-Adder
*
.subckt FULL-ADDER  COUT SOUT CIN XIN YIN

        X_HALF-ADDER1 N$3 SOUT N$220 CIN HALF-ADDER
        X_HALF-ADDER3 N$2 N$220 XIN YIN HALF-ADDER
        X_OR1 COUT N$2 N$3 OR
.ends FULL-ADDER

*
* Component pathname : $UpdatedFiles/default.group/logic.views/4-Bit-Adder
*
.subckt 4-BIT-ADDER  COUT S0 S1 S2 S3 CIN X0 X1 X2 X3 Y0 Y1 Y2 Y3

        X_FULL-ADDER1 N$440 S0 CIN X0 Y0 FULL-ADDER
        X_FULL-ADDER5 COUT S3 N$428 X3 Y3 FULL-ADDER
        X_FULL-ADDER6 N$428 S2 N$433 X2 Y2 FULL-ADDER
        X_FULL-ADDER7 N$433 S1 N$440 X1 Y1 FULL-ADDER
.ends 4-BIT-ADDER

*
* MAIN CELL: Component pathname : $UpdatedFiles/default.group/logic.views/Test_Schematic
*
        V8 N$212 GROUND PATTERN 5 0 0 1n 1n 50n 11111101010
        V7 N$207 GROUND PATTERN 5 0 0 1n 1n 50n 00000101010
        V6 N$211 GROUND PATTERN 5 0 0 1n 1n 50n 01010111101
        V5 N$205 GROUND PATTERN 5 0 0 1n 1n 50n 01010000101
        V4 N$210 GROUND PATTERN 5 0 0 1n 1n 50n 11010010110
        V3 N$213 GROUND PATTERN 5 0 0 1n 1n 50n 01011010010
        V2 N$209 GROUND PATTERN 5 0 0 1n 1n 50n 01100110011
        V1 N$202 GROUND PATTERN 5 0 0 1n 1n 50n 00110011001
        V9 VDD GROUND DC 3.3V
        X_4-BIT-ADDER1 COUT S0 S1 S2 S3 GROUND N$202 N$213 N$205 N$207 N$209
+ N$210 N$211 N$212 4-BIT-ADDER
*
.end
